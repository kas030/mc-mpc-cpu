module add1(a, x);
	input [4:0] a;
	output [4:0] x;
	assign x = a + 5'b1;
endmodule
